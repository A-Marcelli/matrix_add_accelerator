-- ieee packages ------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--use ieee.std_logic_misc.all;
--use ieee.math_real.all;
--use std.textio.all;


entity matrix_add_accelerator is
	generic(


		 );
  port (


  	);
 
 end entity matrix_add_accelerator;

 

 architecture mat_acc of matrix_add_accelerator is 
 	--constants


 	--subtypes


 	--signals


 	--components

 	begin



 end mat_acc;