-- ieee packages ------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Byte_Busters.all;

entity acc_logic is 
	generic(
		);
	port(
		);
end acc_logic;


architecture logic of acc_logic is



begin



end logic;